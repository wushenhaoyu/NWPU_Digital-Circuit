library verilog;
use verilog.vl_types.all;
entity exa4_1 is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : out    vl_logic
    );
end exa4_1;
