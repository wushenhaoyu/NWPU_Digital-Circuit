library verilog;
use verilog.vl_types.all;
entity v5_1_vlg_vec_tst is
end v5_1_vlg_vec_tst;
