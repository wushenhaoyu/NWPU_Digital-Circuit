LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY exa4_1 IS
PORT(A,B:IN STD_LOGIC;
C:OUT STD_LOGIC);
END exa4_1;
ARCHITECTURE fwm OF exa4_1 is
BEGIN 
C<=(NOT A AND B)or(NOT B AND A);
END;