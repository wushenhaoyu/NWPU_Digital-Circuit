library verilog;
use verilog.vl_types.all;
entity \3_3\ is
    port(
        D               : out    vl_logic;
        a               : in     vl_logic;
        b               : in     vl_logic;
        bin             : in     vl_logic;
        \1\             : in     vl_logic;
        \2\             : in     vl_logic;
        \8\             : in     vl_logic;
        \4\             : in     vl_logic;
        Bout            : out    vl_logic
    );
end \3_3\;
