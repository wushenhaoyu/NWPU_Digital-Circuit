library verilog;
use verilog.vl_types.all;
entity \3_2\ is
    port(
        \0\             : out    vl_logic;
        \01\            : in     vl_logic;
        stop            : in     vl_logic;
        \1\             : out    vl_logic;
        \2\             : out    vl_logic;
        \3\             : out    vl_logic;
        \4\             : out    vl_logic;
        \5\             : out    vl_logic;
        \6\             : out    vl_logic;
        Clk             : in     vl_logic
    );
end \3_2\;
