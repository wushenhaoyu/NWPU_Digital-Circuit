library verilog;
use verilog.vl_types.all;
entity exa4_3_vlg_vec_tst is
end exa4_3_vlg_vec_tst;
