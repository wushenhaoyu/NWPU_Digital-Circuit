library verilog;
use verilog.vl_types.all;
entity exa4_1_vlg_check_tst is
    port(
        C               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end exa4_1_vlg_check_tst;
